// nothing yet! :-)